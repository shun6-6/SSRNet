`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/10/18 14:27:27
// Design Name: 
// Module Name: mac_table
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mac_table(
    input           i_clk           ,
    input           i_rst           ,

    input  [47:0]   i_check_mac     , 
    input  [3 :0]   i_check_id      ,
    input           i_check_valid   , 

    output [3 :0]   o_outport       ,
    output          o_result_valid  ,
    output [3 :0]   o_check_id      
);
/******************************function*****************************/

/******************************parameter****************************/

/******************************machine******************************/

/******************************reg**********************************/

/******************************wire*********************************/

/******************************assign*******************************/

/******************************component****************************/

/******************************always*******************************/



endmodule
